module bcd7seg (
	input [7:0] b,
	output reg [13:0] h
);
	assign h[13]=(~b[7]&~b[6]&~b[5]&~b[4])|(~b[7]&~b[6]&~b[5]&b[4])|(~b[7]&b[6]&b[5]&b[4])|(b[7]&b[6]&~b[5]&~b[4]);
	assign h[12]=(~b[7]&~b[6]&~b[5]&b[4])|(~b[7]&~b[6]&b[5]&~b[4])|(~b[7]&~b[6]&b[5]&b[4])|(~b[7]&b[6]&b[5]&b[4])|(b[7]&b[6]&~b[5]&b[4]);
	assign h[11]=(~b[7]&~b[6]&~b[5]&b[4])|(~b[7]&~b[6]&b[5]&b[4])|(~b[7]&b[6]&~b[5]&~b[4])|(~b[7]&b[6]&~b[5]&b[4])|(~b[7]&b[6]&b[5]&b[4])|(b[7]&~b[6]&~b[5]&b[4]);
	assign h[10]=(~b[7]&~b[6]&~b[5]&b[4])|(~b[7]&b[6]&~b[5]&~b[4])|(~b[7]&b[6]&b[5]&b[4])|(b[7]&~b[6]&~b[5]&b[4])|(b[7]&~b[6]&b[5]&~b[4])|(b[7]&b[6]&b[5]&b[4]);
	assign h[9]=(~b[7]&~b[6]&b[5]&~b[4])|(b[7]&b[6]&~b[5]&~b[4])|(b[7]&b[6]&b[5]&~b[4])|(b[7]&b[6]&b[5]&b[4]);
	assign h[8]=(~b[7]&b[6]&~b[5]&b[4])|(~b[7]&b[6]&b[5]&~b[4])|(b[7]&~b[6]&b[5]&b[4])|(b[7]&b[6]&~b[5]&~b[4])|(b[7]&b[6]&b[5]&~b[4])|(b[7]&b[6]&b[5]&b[4]);
	assign h[7]=(~b[7]&~b[6]&~b[5]&b[4])|(~b[7]&b[6]&~b[5]&~b[4])|(b[7]&~b[6]&b[5]&b[4])|(b[7]&b[6]&~b[5]&b[4]);
	assign h[6]=(~b[3]&~b[2]&~b[1]&~b[0])|(~b[3]&~b[2]&~b[1]&b[0])|(~b[3]&b[2]&b[1]&b[0])|(b[3]&b[2]&~b[1]&~b[0]);
	assign h[5]=(~b[3]&~b[2]&~b[1]&b[0])|(~b[3]&~b[2]&b[1]&~b[0])|(~b[3]&~b[2]&b[1]&b[0])|(~b[3]&b[2]&b[1]&b[0])|(b[3]&b[2]&~b[1]&b[0]);
	assign h[4]=(~b[3]&~b[2]&~b[1]&b[0])|(~b[3]&~b[2]&b[1]&b[0])|(~b[3]&b[2]&~b[1]&~b[0])|(~b[3]&b[2]&~b[1]&b[0])|(~b[3]&b[2]&b[1]&b[0])|(b[3]&~b[2]&~b[1]&b[0]);
	assign h[3]=(~b[3]&~b[2]&~b[1]&b[0])|(~b[3]&b[2]&~b[1]&~b[0])|(~b[3]&b[2]&b[1]&b[0])|(b[3]&~b[2]&~b[1]&b[0])|(b[3]&~b[2]&b[1]&~b[0])|(b[3]&b[2]&b[1]&b[0]);
	assign h[2]=(~b[3]&~b[2]&b[1]&~b[0])|(b[3]&b[2]&~b[1]&~b[0])|(b[3]&b[2]&b[1]&~b[0])|(b[3]&b[2]&b[1]&b[0]);
	assign h[1]=(~b[3]&b[2]&~b[1]&b[0])|(~b[3]&b[2]&b[1]&~b[0])|(b[3]&~b[2]&b[1]&b[0])|(b[3]&b[2]&~b[1]&~b[0])|(b[3]&b[2]&b[1]&~b[0])|(b[3]&b[2]&b[1]&b[0]);
	assign h[0]=(~b[3]&~b[2]&~b[1]&b[0])|(~b[3]&b[2]&~b[1]&~b[0])|(b[3]&~b[2]&b[1]&b[0])|(b[3]&b[2]&~b[1]&b[0]);

endmodule

